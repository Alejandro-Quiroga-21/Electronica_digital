`default_nettype none
`define DUMPSTR(x) `"x.vcd`"
`timescale 100ns / 10ns

module Eje_01_tb();

parameter DURATION = 10;


reg clk=0;
always #0.5 clk = ~clk;

// Entradas
reg A_test, B_test;
//Salidas
wire X_test;

Eje_01 UUT (
    .A(A_test),
    .B(B_test),
    .X(X_test)
);

integer  i;
 

initial begin
    // Inicializa las señales
    $dumpfile(`DUMPSTR(`VCD_OUTPUT));
    $dumpvars(0, Eje_01_tb);

    for (i=0;i<4;i=i+1)
        begin
            A_test = i[1];
            B_test = i[0];
            #1;
        end
    //$display ("Current loop # %0d",i);
    A_test = 1'b0;
    B_test = 1'b0;
    #1;
    A_test = 1'b1;
    B_test = 1'b0;
    #1;
    A_test = 1'b1;
    B_test = 1'b1;
    #1;
    A_test = 1'b1;
    B_test = 1'b0;
    #1;
    A_test = 1'b0;
    B_test = 1'b0;
    #1;

    
    
        // Finaliza la simulación
        // $display("Simulación completada.");
    #(DURATION) $display("End of simulation");
    $finish;
    end
    
endmodule