module Eje_01(
    input wire A,B,
    output wire X
);

assign X = A&B;

endmodule